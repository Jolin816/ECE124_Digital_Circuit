library ieee;
use ieee.std_logic_1164.all;

entity seg7_mux is 
port (
	in_1, in_2									: in std_logic_vector (3 downto 0);
	hex_out                             : out std_logic_vector (3 downto 0)
);

end seg7_mux;

architecture  seg7_mux of seg7_mux is

begin

				  
end seg7_mux;
